{"bonuses":[{"Uid":"death","Position":{"X":0.0,"Y":-1.5,"Z":-2.5},"IsEnabled":true},{"Uid":"speedOn","Position":{"X":6.960000038146973,"Y":0.03999999910593033,"Z":2.619999885559082},"IsEnabled":true},{"Uid":"speedOn","Position":{"X":5.0,"Y":-0.004999999888241291,"Z":-6.75},"IsEnabled":true},{"Uid":"point","Position":{"X":-12.0,"Y":0.5,"Z":13.0},"IsEnabled":true},{"Uid":"point","Position":{"X":-2.0,"Y":0.5,"Z":-13.75},"IsEnabled":true},{"Uid":"point","Position":{"X":9.0,"Y":0.5,"Z":13.0},"IsEnabled":true}]}